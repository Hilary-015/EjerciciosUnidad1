----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:31:08 05/15/2022 
-- Design Name: 
-- Module Name:    Promedio - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


--Hilary Calva
entity Promedio is
    Port ( A : in  STD_LOGIC_VECTOR (0 to 3);
           B : in  STD_LOGIC_VECTOR (0 to 3);
           C : out  STD_LOGIC_VECTOR (0 to 3));
end Promedio;

architecture Behavioral of Promedio is

begin


end Behavioral;

