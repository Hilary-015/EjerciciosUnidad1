----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:26:04 05/15/2022 
-- Design Name: 
-- Module Name:    circuito1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


--Hilary Calva

entity circuito1 is
    Port ( A, B : in  STD_LOGIC;
           C : out  STD_LOGIC);
end circuito1;

architecture Behavioral of circuito1 is

begin


end Behavioral;

