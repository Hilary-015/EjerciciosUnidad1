----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:44:27 05/15/2022 
-- Design Name: 
-- Module Name:    MUXVectores - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--Hilary Calva
entity MUXVectores is
    Port ( E : in  STD_LOGIC_VECTOR (0 to 3);
           S : in  STD_LOGIC_VECTOR (0 to 1);
           F : out  STD_LOGIC);
end MUXVectores;

architecture Behavioral of MUXVectores is

begin


end Behavioral;

