----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:50:28 05/15/2022 
-- Design Name: 
-- Module Name:    flujo - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


--Hilary Calva
entity flujo is
    Port ( a0, b0, a1, b1, a2, b2, a3, b3 : in  STD_LOGIC;
           F : out  STD_LOGIC);
end flujo;

architecture Behavioral of flujo is

begin


end Behavioral;

