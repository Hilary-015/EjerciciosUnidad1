----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:28:33 05/15/2022 
-- Design Name: 
-- Module Name:    Proyecto - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--Hilary Calva
entity Proyecto is
    Port ( P0, P1, P2 : in  STD_LOGIC;
           A0, A1 : out  STD_LOGIC;
           X : inout  STD_LOGIC);
end Proyecto;

architecture Behavioral of Proyecto is

begin


end Behavioral;

